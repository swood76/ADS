-- nios.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity nios is
	port (
		clk_clk                           : in  std_logic := '0'; --                        clk.clk
		led_external_connection_export    : out std_logic;        --    led_external_connection.export
		reset_reset_n                     : in  std_logic := '0'; --                      reset.reset_n
		switch_external_connection_export : in  std_logic := '0'  -- switch_external_connection.export
	);
end entity nios;

architecture rtl of nios is
	component nios_led is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic                                         -- export
		);
	end component nios_led;

	component nios_nios2e is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(14 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(14 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component nios_nios2e;

	component nios_onchip_memory is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(11 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component nios_onchip_memory;

	component nios_switch is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic                     := 'X'              -- export
		);
	end component nios_switch;

	component nios_uart is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component nios_uart;

	component nios_mm_interconnect_0 is
		port (
			clk_0_clk_clk                            : in  std_logic                     := 'X';             -- clk
			nios2e_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			nios2e_data_master_address               : in  std_logic_vector(14 downto 0) := (others => 'X'); -- address
			nios2e_data_master_waitrequest           : out std_logic;                                        -- waitrequest
			nios2e_data_master_byteenable            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			nios2e_data_master_read                  : in  std_logic                     := 'X';             -- read
			nios2e_data_master_readdata              : out std_logic_vector(31 downto 0);                    -- readdata
			nios2e_data_master_write                 : in  std_logic                     := 'X';             -- write
			nios2e_data_master_writedata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			nios2e_data_master_debugaccess           : in  std_logic                     := 'X';             -- debugaccess
			nios2e_instruction_master_address        : in  std_logic_vector(14 downto 0) := (others => 'X'); -- address
			nios2e_instruction_master_waitrequest    : out std_logic;                                        -- waitrequest
			nios2e_instruction_master_read           : in  std_logic                     := 'X';             -- read
			nios2e_instruction_master_readdata       : out std_logic_vector(31 downto 0);                    -- readdata
			led_s1_address                           : out std_logic_vector(1 downto 0);                     -- address
			led_s1_write                             : out std_logic;                                        -- write
			led_s1_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			led_s1_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			led_s1_chipselect                        : out std_logic;                                        -- chipselect
			nios2e_debug_mem_slave_address           : out std_logic_vector(8 downto 0);                     -- address
			nios2e_debug_mem_slave_write             : out std_logic;                                        -- write
			nios2e_debug_mem_slave_read              : out std_logic;                                        -- read
			nios2e_debug_mem_slave_readdata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nios2e_debug_mem_slave_writedata         : out std_logic_vector(31 downto 0);                    -- writedata
			nios2e_debug_mem_slave_byteenable        : out std_logic_vector(3 downto 0);                     -- byteenable
			nios2e_debug_mem_slave_waitrequest       : in  std_logic                     := 'X';             -- waitrequest
			nios2e_debug_mem_slave_debugaccess       : out std_logic;                                        -- debugaccess
			onchip_memory_s1_address                 : out std_logic_vector(11 downto 0);                    -- address
			onchip_memory_s1_write                   : out std_logic;                                        -- write
			onchip_memory_s1_readdata                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_memory_s1_writedata               : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_memory_s1_byteenable              : out std_logic_vector(3 downto 0);                     -- byteenable
			onchip_memory_s1_chipselect              : out std_logic;                                        -- chipselect
			onchip_memory_s1_clken                   : out std_logic;                                        -- clken
			switch_s1_address                        : out std_logic_vector(1 downto 0);                     -- address
			switch_s1_readdata                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			uart_avalon_jtag_slave_address           : out std_logic_vector(0 downto 0);                     -- address
			uart_avalon_jtag_slave_write             : out std_logic;                                        -- write
			uart_avalon_jtag_slave_read              : out std_logic;                                        -- read
			uart_avalon_jtag_slave_readdata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			uart_avalon_jtag_slave_writedata         : out std_logic_vector(31 downto 0);                    -- writedata
			uart_avalon_jtag_slave_waitrequest       : in  std_logic                     := 'X';             -- waitrequest
			uart_avalon_jtag_slave_chipselect        : out std_logic                                         -- chipselect
		);
	end component nios_mm_interconnect_0;

	component nios_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component nios_irq_mapper;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal nios2e_data_master_readdata                              : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2e_data_master_readdata -> nios2e:d_readdata
	signal nios2e_data_master_waitrequest                           : std_logic;                     -- mm_interconnect_0:nios2e_data_master_waitrequest -> nios2e:d_waitrequest
	signal nios2e_data_master_debugaccess                           : std_logic;                     -- nios2e:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2e_data_master_debugaccess
	signal nios2e_data_master_address                               : std_logic_vector(14 downto 0); -- nios2e:d_address -> mm_interconnect_0:nios2e_data_master_address
	signal nios2e_data_master_byteenable                            : std_logic_vector(3 downto 0);  -- nios2e:d_byteenable -> mm_interconnect_0:nios2e_data_master_byteenable
	signal nios2e_data_master_read                                  : std_logic;                     -- nios2e:d_read -> mm_interconnect_0:nios2e_data_master_read
	signal nios2e_data_master_write                                 : std_logic;                     -- nios2e:d_write -> mm_interconnect_0:nios2e_data_master_write
	signal nios2e_data_master_writedata                             : std_logic_vector(31 downto 0); -- nios2e:d_writedata -> mm_interconnect_0:nios2e_data_master_writedata
	signal nios2e_instruction_master_readdata                       : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2e_instruction_master_readdata -> nios2e:i_readdata
	signal nios2e_instruction_master_waitrequest                    : std_logic;                     -- mm_interconnect_0:nios2e_instruction_master_waitrequest -> nios2e:i_waitrequest
	signal nios2e_instruction_master_address                        : std_logic_vector(14 downto 0); -- nios2e:i_address -> mm_interconnect_0:nios2e_instruction_master_address
	signal nios2e_instruction_master_read                           : std_logic;                     -- nios2e:i_read -> mm_interconnect_0:nios2e_instruction_master_read
	signal mm_interconnect_0_nios2e_debug_mem_slave_readdata        : std_logic_vector(31 downto 0); -- nios2e:debug_mem_slave_readdata -> mm_interconnect_0:nios2e_debug_mem_slave_readdata
	signal mm_interconnect_0_nios2e_debug_mem_slave_waitrequest     : std_logic;                     -- nios2e:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2e_debug_mem_slave_waitrequest
	signal mm_interconnect_0_nios2e_debug_mem_slave_debugaccess     : std_logic;                     -- mm_interconnect_0:nios2e_debug_mem_slave_debugaccess -> nios2e:debug_mem_slave_debugaccess
	signal mm_interconnect_0_nios2e_debug_mem_slave_address         : std_logic_vector(8 downto 0);  -- mm_interconnect_0:nios2e_debug_mem_slave_address -> nios2e:debug_mem_slave_address
	signal mm_interconnect_0_nios2e_debug_mem_slave_read            : std_logic;                     -- mm_interconnect_0:nios2e_debug_mem_slave_read -> nios2e:debug_mem_slave_read
	signal mm_interconnect_0_nios2e_debug_mem_slave_byteenable      : std_logic_vector(3 downto 0);  -- mm_interconnect_0:nios2e_debug_mem_slave_byteenable -> nios2e:debug_mem_slave_byteenable
	signal mm_interconnect_0_nios2e_debug_mem_slave_write           : std_logic;                     -- mm_interconnect_0:nios2e_debug_mem_slave_write -> nios2e:debug_mem_slave_write
	signal mm_interconnect_0_nios2e_debug_mem_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2e_debug_mem_slave_writedata -> nios2e:debug_mem_slave_writedata
	signal mm_interconnect_0_uart_avalon_jtag_slave_chipselect      : std_logic;                     -- mm_interconnect_0:uart_avalon_jtag_slave_chipselect -> uart:av_chipselect
	signal mm_interconnect_0_uart_avalon_jtag_slave_readdata        : std_logic_vector(31 downto 0); -- uart:av_readdata -> mm_interconnect_0:uart_avalon_jtag_slave_readdata
	signal mm_interconnect_0_uart_avalon_jtag_slave_waitrequest     : std_logic;                     -- uart:av_waitrequest -> mm_interconnect_0:uart_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_uart_avalon_jtag_slave_address         : std_logic_vector(0 downto 0);  -- mm_interconnect_0:uart_avalon_jtag_slave_address -> uart:av_address
	signal mm_interconnect_0_uart_avalon_jtag_slave_read            : std_logic;                     -- mm_interconnect_0:uart_avalon_jtag_slave_read -> mm_interconnect_0_uart_avalon_jtag_slave_read:in
	signal mm_interconnect_0_uart_avalon_jtag_slave_write           : std_logic;                     -- mm_interconnect_0:uart_avalon_jtag_slave_write -> mm_interconnect_0_uart_avalon_jtag_slave_write:in
	signal mm_interconnect_0_uart_avalon_jtag_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:uart_avalon_jtag_slave_writedata -> uart:av_writedata
	signal mm_interconnect_0_onchip_memory_s1_chipselect            : std_logic;                     -- mm_interconnect_0:onchip_memory_s1_chipselect -> onchip_memory:chipselect
	signal mm_interconnect_0_onchip_memory_s1_readdata              : std_logic_vector(31 downto 0); -- onchip_memory:readdata -> mm_interconnect_0:onchip_memory_s1_readdata
	signal mm_interconnect_0_onchip_memory_s1_address               : std_logic_vector(11 downto 0); -- mm_interconnect_0:onchip_memory_s1_address -> onchip_memory:address
	signal mm_interconnect_0_onchip_memory_s1_byteenable            : std_logic_vector(3 downto 0);  -- mm_interconnect_0:onchip_memory_s1_byteenable -> onchip_memory:byteenable
	signal mm_interconnect_0_onchip_memory_s1_write                 : std_logic;                     -- mm_interconnect_0:onchip_memory_s1_write -> onchip_memory:write
	signal mm_interconnect_0_onchip_memory_s1_writedata             : std_logic_vector(31 downto 0); -- mm_interconnect_0:onchip_memory_s1_writedata -> onchip_memory:writedata
	signal mm_interconnect_0_onchip_memory_s1_clken                 : std_logic;                     -- mm_interconnect_0:onchip_memory_s1_clken -> onchip_memory:clken
	signal mm_interconnect_0_led_s1_chipselect                      : std_logic;                     -- mm_interconnect_0:led_s1_chipselect -> led:chipselect
	signal mm_interconnect_0_led_s1_readdata                        : std_logic_vector(31 downto 0); -- led:readdata -> mm_interconnect_0:led_s1_readdata
	signal mm_interconnect_0_led_s1_address                         : std_logic_vector(1 downto 0);  -- mm_interconnect_0:led_s1_address -> led:address
	signal mm_interconnect_0_led_s1_write                           : std_logic;                     -- mm_interconnect_0:led_s1_write -> mm_interconnect_0_led_s1_write:in
	signal mm_interconnect_0_led_s1_writedata                       : std_logic_vector(31 downto 0); -- mm_interconnect_0:led_s1_writedata -> led:writedata
	signal mm_interconnect_0_switch_s1_readdata                     : std_logic_vector(31 downto 0); -- switch:readdata -> mm_interconnect_0:switch_s1_readdata
	signal mm_interconnect_0_switch_s1_address                      : std_logic_vector(1 downto 0);  -- mm_interconnect_0:switch_s1_address -> switch:address
	signal irq_mapper_receiver0_irq                                 : std_logic;                     -- uart:av_irq -> irq_mapper:receiver0_irq
	signal nios2e_irq_irq                                           : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> nios2e:irq
	signal rst_controller_reset_out_reset                           : std_logic;                     -- rst_controller:reset_out -> [irq_mapper:reset, mm_interconnect_0:nios2e_reset_reset_bridge_in_reset_reset, onchip_memory:reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                       : std_logic;                     -- rst_controller:reset_req -> [nios2e:reset_req, onchip_memory:reset_req, rst_translator:reset_req_in]
	signal reset_reset_n_ports_inv                                  : std_logic;                     -- reset_reset_n:inv -> rst_controller:reset_in0
	signal mm_interconnect_0_uart_avalon_jtag_slave_read_ports_inv  : std_logic;                     -- mm_interconnect_0_uart_avalon_jtag_slave_read:inv -> uart:av_read_n
	signal mm_interconnect_0_uart_avalon_jtag_slave_write_ports_inv : std_logic;                     -- mm_interconnect_0_uart_avalon_jtag_slave_write:inv -> uart:av_write_n
	signal mm_interconnect_0_led_s1_write_ports_inv                 : std_logic;                     -- mm_interconnect_0_led_s1_write:inv -> led:write_n
	signal rst_controller_reset_out_reset_ports_inv                 : std_logic;                     -- rst_controller_reset_out_reset:inv -> [led:reset_n, nios2e:reset_n, switch:reset_n, uart:rst_n]

begin

	led : component nios_led
		port map (
			clk        => clk_clk,                                  --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_0_led_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_led_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_led_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_led_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_led_s1_readdata,        --                    .readdata
			out_port   => led_external_connection_export            -- external_connection.export
		);

	nios2e : component nios_nios2e
		port map (
			clk                                 => clk_clk,                                              --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,             --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                   --                          .reset_req
			d_address                           => nios2e_data_master_address,                           --               data_master.address
			d_byteenable                        => nios2e_data_master_byteenable,                        --                          .byteenable
			d_read                              => nios2e_data_master_read,                              --                          .read
			d_readdata                          => nios2e_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => nios2e_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => nios2e_data_master_write,                             --                          .write
			d_writedata                         => nios2e_data_master_writedata,                         --                          .writedata
			debug_mem_slave_debugaccess_to_roms => nios2e_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => nios2e_instruction_master_address,                    --        instruction_master.address
			i_read                              => nios2e_instruction_master_read,                       --                          .read
			i_readdata                          => nios2e_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => nios2e_instruction_master_waitrequest,                --                          .waitrequest
			irq                                 => nios2e_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => open,                                                 --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_nios2e_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_nios2e_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_nios2e_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_nios2e_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_nios2e_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_nios2e_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_nios2e_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_nios2e_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                  -- custom_instruction_master.readra
		);

	onchip_memory : component nios_onchip_memory
		port map (
			clk        => clk_clk,                                       --   clk1.clk
			address    => mm_interconnect_0_onchip_memory_s1_address,    --     s1.address
			clken      => mm_interconnect_0_onchip_memory_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_onchip_memory_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_onchip_memory_s1_write,      --       .write
			readdata   => mm_interconnect_0_onchip_memory_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_onchip_memory_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_onchip_memory_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,                -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req,            --       .reset_req
			freeze     => '0'                                            -- (terminated)
		);

	switch : component nios_switch
		port map (
			clk      => clk_clk,                                  --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_switch_s1_address,      --                  s1.address
			readdata => mm_interconnect_0_switch_s1_readdata,     --                    .readdata
			in_port  => switch_external_connection_export         -- external_connection.export
		);

	uart : component nios_uart
		port map (
			clk            => clk_clk,                                                  --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                 --             reset.reset_n
			av_chipselect  => mm_interconnect_0_uart_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_uart_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_uart_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_uart_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_uart_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_uart_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_uart_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver0_irq                                  --               irq.irq
		);

	mm_interconnect_0 : component nios_mm_interconnect_0
		port map (
			clk_0_clk_clk                            => clk_clk,                                              --                          clk_0_clk.clk
			nios2e_reset_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                       -- nios2e_reset_reset_bridge_in_reset.reset
			nios2e_data_master_address               => nios2e_data_master_address,                           --                 nios2e_data_master.address
			nios2e_data_master_waitrequest           => nios2e_data_master_waitrequest,                       --                                   .waitrequest
			nios2e_data_master_byteenable            => nios2e_data_master_byteenable,                        --                                   .byteenable
			nios2e_data_master_read                  => nios2e_data_master_read,                              --                                   .read
			nios2e_data_master_readdata              => nios2e_data_master_readdata,                          --                                   .readdata
			nios2e_data_master_write                 => nios2e_data_master_write,                             --                                   .write
			nios2e_data_master_writedata             => nios2e_data_master_writedata,                         --                                   .writedata
			nios2e_data_master_debugaccess           => nios2e_data_master_debugaccess,                       --                                   .debugaccess
			nios2e_instruction_master_address        => nios2e_instruction_master_address,                    --          nios2e_instruction_master.address
			nios2e_instruction_master_waitrequest    => nios2e_instruction_master_waitrequest,                --                                   .waitrequest
			nios2e_instruction_master_read           => nios2e_instruction_master_read,                       --                                   .read
			nios2e_instruction_master_readdata       => nios2e_instruction_master_readdata,                   --                                   .readdata
			led_s1_address                           => mm_interconnect_0_led_s1_address,                     --                             led_s1.address
			led_s1_write                             => mm_interconnect_0_led_s1_write,                       --                                   .write
			led_s1_readdata                          => mm_interconnect_0_led_s1_readdata,                    --                                   .readdata
			led_s1_writedata                         => mm_interconnect_0_led_s1_writedata,                   --                                   .writedata
			led_s1_chipselect                        => mm_interconnect_0_led_s1_chipselect,                  --                                   .chipselect
			nios2e_debug_mem_slave_address           => mm_interconnect_0_nios2e_debug_mem_slave_address,     --             nios2e_debug_mem_slave.address
			nios2e_debug_mem_slave_write             => mm_interconnect_0_nios2e_debug_mem_slave_write,       --                                   .write
			nios2e_debug_mem_slave_read              => mm_interconnect_0_nios2e_debug_mem_slave_read,        --                                   .read
			nios2e_debug_mem_slave_readdata          => mm_interconnect_0_nios2e_debug_mem_slave_readdata,    --                                   .readdata
			nios2e_debug_mem_slave_writedata         => mm_interconnect_0_nios2e_debug_mem_slave_writedata,   --                                   .writedata
			nios2e_debug_mem_slave_byteenable        => mm_interconnect_0_nios2e_debug_mem_slave_byteenable,  --                                   .byteenable
			nios2e_debug_mem_slave_waitrequest       => mm_interconnect_0_nios2e_debug_mem_slave_waitrequest, --                                   .waitrequest
			nios2e_debug_mem_slave_debugaccess       => mm_interconnect_0_nios2e_debug_mem_slave_debugaccess, --                                   .debugaccess
			onchip_memory_s1_address                 => mm_interconnect_0_onchip_memory_s1_address,           --                   onchip_memory_s1.address
			onchip_memory_s1_write                   => mm_interconnect_0_onchip_memory_s1_write,             --                                   .write
			onchip_memory_s1_readdata                => mm_interconnect_0_onchip_memory_s1_readdata,          --                                   .readdata
			onchip_memory_s1_writedata               => mm_interconnect_0_onchip_memory_s1_writedata,         --                                   .writedata
			onchip_memory_s1_byteenable              => mm_interconnect_0_onchip_memory_s1_byteenable,        --                                   .byteenable
			onchip_memory_s1_chipselect              => mm_interconnect_0_onchip_memory_s1_chipselect,        --                                   .chipselect
			onchip_memory_s1_clken                   => mm_interconnect_0_onchip_memory_s1_clken,             --                                   .clken
			switch_s1_address                        => mm_interconnect_0_switch_s1_address,                  --                          switch_s1.address
			switch_s1_readdata                       => mm_interconnect_0_switch_s1_readdata,                 --                                   .readdata
			uart_avalon_jtag_slave_address           => mm_interconnect_0_uart_avalon_jtag_slave_address,     --             uart_avalon_jtag_slave.address
			uart_avalon_jtag_slave_write             => mm_interconnect_0_uart_avalon_jtag_slave_write,       --                                   .write
			uart_avalon_jtag_slave_read              => mm_interconnect_0_uart_avalon_jtag_slave_read,        --                                   .read
			uart_avalon_jtag_slave_readdata          => mm_interconnect_0_uart_avalon_jtag_slave_readdata,    --                                   .readdata
			uart_avalon_jtag_slave_writedata         => mm_interconnect_0_uart_avalon_jtag_slave_writedata,   --                                   .writedata
			uart_avalon_jtag_slave_waitrequest       => mm_interconnect_0_uart_avalon_jtag_slave_waitrequest, --                                   .waitrequest
			uart_avalon_jtag_slave_chipselect        => mm_interconnect_0_uart_avalon_jtag_slave_chipselect   --                                   .chipselect
		);

	irq_mapper : component nios_irq_mapper
		port map (
			clk           => clk_clk,                        --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			sender_irq    => nios2e_irq_irq                  --    sender.irq
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_uart_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_uart_avalon_jtag_slave_read;

	mm_interconnect_0_uart_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_uart_avalon_jtag_slave_write;

	mm_interconnect_0_led_s1_write_ports_inv <= not mm_interconnect_0_led_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of nios
